// tb/tb_cpu.sv
`timescale 1ns/1ps

module tb_cpu;
  //-------------------------------------------------------------------------
  // Clock & reset
  //-------------------------------------------------------------------------
  logic clk   = 0;
  logic reset = 1;

  always #5 clk = ~clk;  // 100 MHz

  initial begin
    #20 reset = 0;       // release reset after 20 ns
  end

  //-------------------------------------------------------------------------
  // DUT instantiation
  //-------------------------------------------------------------------------
  cpu dut (
    .clk   (clk),
    .reset (reset)
  );

  //-------------------------------------------------------------------------
  // Waveform dumping
  //-------------------------------------------------------------------------
  initial begin
    $dumpfile("tb_cpu.vcd");
    $dumpvars(0, tb_cpu);
  end

  //-------------------------------------------------------------------------
  // Test timeout / finish
  //-------------------------------------------------------------------------
  initial begin
    #10000;
    $display("**** TIMEOUT ****");
    $finish;
  end
endmodule
